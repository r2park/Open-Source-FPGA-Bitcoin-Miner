library verilog;
use verilog.vl_types.all;
entity test_fpgaminer_top is
end test_fpgaminer_top;
